`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:53:07 11/29/2020 
// Design Name: 
// Module Name:    MFCMP1D 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MFCMP1D(
	input [3:0] mfcmp1dSel,
	input [31:0] V1,
	input [31:0] ALUC_M,
	input [31:0] pc4_M,
	input [31:0] ALUC_W,
	input [31:0] DMRD_W,
	output [31:0] mfcmp1d
    );


endmodule
